CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
10 0 10 150 10
170 80 1438 831
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
338 176 451 273
42991634 0
0
6 Title:
5 Name:
0
0
0
31
13 Logic Switch~
5 68 455 0 1 11
0 16
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3277 0 0
2
45449.4 0
0
13 Logic Switch~
5 86 268 0 1 11
0 20
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4212 0 0
2
45449.4 1
0
13 Logic Switch~
5 88 122 0 10 11
0 21 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
4720 0 0
2
45449.4 2
0
14 Logic Display~
6 701 979 0 1 2
10 2
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L12
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5551 0 0
2
5.90126e-315 0
0
14 Logic Display~
6 587 979 0 1 2
10 3
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L11
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6986 0 0
2
5.90126e-315 5.26354e-315
0
14 Logic Display~
6 455 981 0 1 2
10 4
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L10
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8745 0 0
2
5.90126e-315 5.30499e-315
0
14 Logic Display~
6 334 985 0 1 2
10 5
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L9
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9592 0 0
2
5.90126e-315 5.32571e-315
0
14 Logic Display~
6 695 901 0 1 2
10 7
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L8
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8748 0 0
2
5.90126e-315 5.34643e-315
0
14 Logic Display~
6 582 903 0 1 2
10 8
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L7
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7168 0 0
2
5.90126e-315 5.3568e-315
0
14 Logic Display~
6 452 905 0 1 2
10 9
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
631 0 0
2
5.90126e-315 5.36716e-315
0
14 Logic Display~
6 332 905 0 1 2
10 10
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9466 0 0
2
5.90126e-315 5.37752e-315
0
12 D Flip-Flop~
219 595 825 0 4 9
0 8 6 2 7
0
0 0 4720 0
3 DFF
-10 -53 11 -45
2 U8
-7 -55 7 -47
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
11 typeDigital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 0 1 0 0 0
1 U
3266 0 0
2
5.90126e-315 5.38788e-315
0
12 D Flip-Flop~
219 465 825 0 4 9
0 9 6 3 8
0
0 0 4720 0
3 DFF
-10 -53 11 -45
2 U7
-7 -55 7 -47
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
11 typeDigital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 0 1 0 0 0
1 U
7693 0 0
2
5.90126e-315 5.39306e-315
0
12 D Flip-Flop~
219 344 825 0 4 9
0 10 6 4 9
0
0 0 4720 0
3 DFF
-10 -53 11 -45
2 U6
-7 -55 7 -47
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
11 typeDigital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 0 1 0 0 0
1 U
3723 0 0
2
5.90126e-315 5.39824e-315
0
12 D Flip-Flop~
219 232 825 0 4 9
0 2 6 5 10
0
0 0 4720 0
3 DFF
-10 -53 11 -45
2 U5
-7 -55 7 -47
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
11 typeDigital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 0 1 0 0 0
1 U
3440 0 0
2
5.90126e-315 5.40342e-315
0
7 Pulser~
4 50 816 0 10 12
0 25 26 6 27 0 0 20 20 13
7
0
0 0 4656 0
0
3 V10
-11 -28 10 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
6263 0 0
2
45449.4 3
0
14 Logic Display~
6 631 564 0 1 2
10 12
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4900 0 0
2
45449.4 4
0
14 Logic Display~
6 620 422 0 1 2
10 11
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8783 0 0
2
45449.4 5
0
10 2-In NAND~
219 472 587 0 3 22
0 11 14 12
0
0 0 624 0
6 74LS00
-14 -24 28 -16
3 U4D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 4 0
1 U
3221 0 0
2
45449.4 6
0
10 2-In NAND~
219 469 448 0 3 22
0 13 12 11
0
0 0 624 0
6 74LS00
-14 -24 28 -16
3 U4C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 4 0
1 U
3215 0 0
2
45449.4 7
0
10 2-In NAND~
219 304 446 0 3 22
0 16 15 13
0
0 0 624 0
6 74LS00
-14 -24 28 -16
3 U4B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 4 0
1 U
7903 0 0
2
45449.4 8
0
10 2-In NAND~
219 302 584 0 3 22
0 15 17 14
0
0 0 624 0
6 74LS00
-14 -24 28 -16
3 U4A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
7121 0 0
2
45449.4 9
0
9 Inverter~
13 118 592 0 2 22
0 16 17
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U3A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 3 0
1 U
4484 0 0
2
45449.4 10
0
7 Pulser~
4 135 523 0 10 12
0 28 29 15 30 0 0 5 5 3
8
0
0 0 4656 0
0
2 V5
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
5996 0 0
2
45449.4 11
0
14 Logic Display~
6 560 221 0 1 2
10 19
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7804 0 0
2
45449.4 12
0
14 Logic Display~
6 555 118 0 1 2
10 18
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5523 0 0
2
45449.4 13
0
7 Pulser~
4 157 198 0 10 12
0 31 32 22 33 0 0 5 5 3
8
0
0 0 4656 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
3330 0 0
2
45449.4 14
0
9 2-In NOR~
219 404 143 0 3 22
0 23 19 18
0
0 0 624 0
6 74LS02
-21 -24 21 -16
3 U2B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
3465 0 0
2
45449.4 15
0
9 2-In NOR~
219 402 249 0 3 22
0 18 24 19
0
0 0 624 0
6 74LS02
-21 -24 21 -16
3 U2A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 3 2 1 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
8396 0 0
2
45449.4 16
0
9 2-In AND~
219 257 259 0 3 22
0 22 20 24
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U1B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
3685 0 0
2
45449.4 17
0
9 2-In AND~
219 259 135 0 3 22
0 21 22 23
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U1A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
7849 0 0
2
45449.4 18
0
37
0 1 2 0 0 4096 0 0 4 6 0 4
629 807
629 1005
701 1005
701 997
3 1 3 0 0 8320 0 13 5 0 0 5
495 807
505 807
505 1005
587 1005
587 997
3 1 4 0 0 8320 0 14 6 0 0 5
374 807
383 807
383 1007
455 1007
455 999
3 1 5 0 0 8320 0 15 7 0 0 5
262 807
268 807
268 1011
334 1011
334 1003
0 2 6 0 0 4096 0 0 12 12 0 4
433 822
563 822
563 807
571 807
3 1 2 0 0 12416 0 12 15 0 0 6
625 807
629 807
629 755
200 755
200 789
208 789
1 4 7 0 0 12416 0 8 12 0 0 5
695 919
695 923
666 923
666 789
619 789
1 0 8 0 0 12416 0 9 0 0 11 4
582 921
582 925
519 925
519 789
1 0 9 0 0 12416 0 10 0 0 13 4
452 923
452 927
396 927
396 789
1 0 10 0 0 12416 0 11 0 0 15 4
332 923
332 927
281 927
281 789
4 1 8 0 0 0 0 13 12 0 0 2
489 789
571 789
0 2 6 0 0 0 0 0 13 14 0 4
312 822
433 822
433 807
441 807
4 1 9 0 0 0 0 14 13 0 0 2
368 789
441 789
0 2 6 0 0 8320 0 0 14 16 0 5
111 807
111 822
312 822
312 807
320 807
4 1 10 0 0 0 0 15 14 0 0 2
256 789
320 789
2 3 6 0 0 0 0 15 16 0 0 2
208 807
74 807
1 0 11 0 0 12288 0 19 0 0 19 5
448 578
441 578
441 532
546 532
546 448
2 0 12 0 0 12288 0 20 0 0 20 4
445 457
445 490
533 490
533 587
3 1 11 0 0 4224 0 20 18 0 0 3
496 448
620 448
620 440
3 1 12 0 0 4224 0 19 17 0 0 3
499 587
631 587
631 582
3 1 13 0 0 4224 0 21 20 0 0 4
331 446
437 446
437 439
445 439
3 2 14 0 0 4224 0 22 19 0 0 4
329 584
440 584
440 596
448 596
3 2 15 0 0 4224 0 24 21 0 0 4
159 514
270 514
270 455
280 455
3 1 15 0 0 0 0 24 22 0 0 4
159 514
270 514
270 575
278 575
0 1 16 0 0 8320 0 0 21 27 0 3
85 455
85 437
280 437
2 2 17 0 0 4224 0 23 22 0 0 4
139 592
268 592
268 593
278 593
1 1 16 0 0 0 0 1 23 0 0 4
80 455
85 455
85 592
103 592
1 0 18 0 0 12288 0 29 0 0 31 5
389 240
385 240
385 196
473 196
473 143
2 0 19 0 0 12288 0 28 0 0 30 5
391 152
382 152
382 180
452 180
452 249
3 1 19 0 0 4224 0 29 25 0 0 5
441 249
545 249
545 250
560 250
560 239
3 1 18 0 0 4224 0 28 26 0 0 3
443 143
555 143
555 136
1 2 20 0 0 4224 0 2 30 0 0 2
98 268
233 268
1 1 21 0 0 4224 0 3 31 0 0 4
100 122
227 122
227 126
235 126
1 3 22 0 0 8320 0 30 27 0 0 4
233 250
222 250
222 189
181 189
2 3 22 0 0 0 0 31 27 0 0 4
235 144
221 144
221 189
181 189
3 1 23 0 0 12416 0 31 28 0 0 4
280 135
295 135
295 134
391 134
3 2 24 0 0 4224 0 30 29 0 0 4
278 259
352 259
352 258
389 258
15
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
30 756 69 780
37 761 61 777
3 CLK
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 21
7 645 196 669
17 653 185 669
21 REPLICADO DE CIRCUITO
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
612 509 649 533
622 517 638 533
2 Q'
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
605 366 634 390
615 374 623 390
1 Q
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
116 463 161 487
126 471 150 487
3 CLK
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
136 138 181 162
146 146 170 162
3 CLK
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
543 169 580 193
553 177 569 193
2 Q'
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
539 64 568 88
549 72 557 88
1 Q
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 11
13 354 122 378
23 362 111 378
11 FLIP FLOP D
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
58 280 119 304
68 288 108 304
5 RESET
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
65 60 110 84
75 68 99 84
3 SET
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 12
11 7 128 31
21 15 117 31
12 FLIP FLOP RS
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 21
271 689 454 713
278 695 446 711
21 FLIPFLOPS EN PARALELO
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 15
254 712 389 736
261 718 381 734
15 ultimo flipflop
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 13
384 712 503 736
391 717 495 733
13 retroalimenta
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
