CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
1140 80 30 150 10
253 80 1438 831
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
5 4 0.500000 0.500000
253 80 1438 831
42991634 0
0
6 Title:
5 Name:
0
0
0
25
9 CA 7-Seg~
184 1891 127 0 18 19
10 35 34 33 32 31 30 3 79 80
0 0 0 0 0 0 2 2 2
0
0 0 21104 0
7 AMBERCA
9 -41 58 -33
5 DISP6
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
5130 0 0
2
45461.5 0
0
9 2-In AND~
219 475 463 0 3 22
0 7 8 6
0
0 0 624 90
6 74LS08
-21 -24 21 -16
4 U10D
17 -5 45 3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 2 0
1 U
391 0 0
2
45461.5 2
0
8 2-In OR~
219 480 389 0 3 22
0 6 9 5
0
0 0 624 90
6 74LS32
-21 -24 21 -16
4 U15A
29 -3 57 5
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
3124 0 0
2
45461.5 3
0
9 2-In AND~
219 595 384 0 3 22
0 11 10 9
0
0 0 624 270
6 74LS08
-21 -24 21 -16
4 U10C
17 -4 45 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 2 0
1 U
3421 0 0
2
45461.5 4
0
6 74LS47
187 1822 244 0 14 29
0 27 28 26 29 81 82 3 30 31
32 33 34 35 83
0
0 0 4848 0
6 74LS47
-21 -60 21 -52
3 U14
-10 -61 11 -53
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
8157 0 0
2
45461.5 5
0
7 74LS193
137 1707 200 0 14 29
0 2 84 85 14 86 87 88 89 90
91 27 28 26 29
0
0 0 4848 0
7 74LS193
-24 -51 25 -43
3 U13
-10 -52 11 -44
0
15 DVCC=16;DGND=8;
122 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 5 4 11 14 9 10 1 15 12
13 7 6 2 3 5 4 11 14 9
10 1 15 12 13 7 6 2 3 0
65 0 0 512 1 0 0 0
1 U
5572 0 0
2
45461.5 6
0
9 2-In AND~
219 1714 299 0 3 22
0 26 27 14
0
0 0 624 180
6 74LS08
-21 -24 21 -16
4 U10B
-16 -25 12 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
8901 0 0
2
45461.5 7
0
7 74LS193
137 1432 212 0 14 29
0 14 92 93 13 94 95 96 97 98
99 17 16 15 18
0
0 0 4848 0
7 74LS193
-24 -51 25 -43
3 U12
-10 -52 11 -44
0
15 DVCC=16;DGND=8;
122 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 5 4 11 14 9 10 1 15 12
13 7 6 2 3 5 4 11 14 9
10 1 15 12 13 7 6 2 3 0
65 0 0 512 1 0 0 0
1 U
7361 0 0
2
45461.5 8
0
9 CA 7-Seg~
184 1615 145 0 18 19
10 25 24 23 22 21 20 19 100 101
0 0 0 0 0 0 2 2 2
0
0 0 21104 0
7 AMBERCA
9 -41 58 -33
5 DISP5
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
4747 0 0
2
45461.5 9
0
6 74LS47
187 1547 256 0 14 29
0 17 16 15 18 102 103 19 20 21
22 23 24 25 104
0
0 0 4848 0
6 74LS47
-21 -60 21 -52
3 U11
-10 -61 11 -53
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
972 0 0
2
45461.5 10
0
9 2-In AND~
219 1436 310 0 3 22
0 16 15 13
0
0 0 624 180
6 74LS08
-21 -24 21 -16
4 U10A
-16 -25 12 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
3472 0 0
2
45461.5 11
0
6 74LS47
187 657 264 0 14 29
0 11 8 10 46 105 106 47 48 49
50 51 52 53 107
0
0 0 4848 0
6 74LS47
-21 -60 21 -52
2 U9
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
9998 0 0
2
45461.5 12
0
9 CA 7-Seg~
184 725 153 0 18 19
10 53 52 51 50 49 48 47 108 109
0 0 0 0 0 0 2 2 2
0
0 0 21104 0
7 AMBERCA
9 -41 58 -33
5 DISP4
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
3536 0 0
2
45461.5 13
0
7 74LS193
137 542 220 0 14 29
0 4 110 111 5 112 113 114 115 116
117 11 8 10 46
0
0 0 4848 0
7 74LS193
-24 -51 25 -43
2 U8
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
122 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 5 4 11 14 9 10 1 15 12
13 7 6 2 3 5 4 11 14 9
10 1 15 12 13 7 6 2 3 0
65 0 0 512 1 0 0 0
1 U
4597 0 0
2
45461.5 14
0
7 74LS193
137 267 232 0 14 29
0 5 118 119 6 120 121 122 123 124
125 36 37 7 38
0
0 0 4848 0
7 74LS193
-24 -51 25 -43
2 U7
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
122 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 5 4 11 14 9 10 1 15 12
13 7 6 2 3 5 4 11 14 9
10 1 15 12 13 7 6 2 3 0
65 0 0 512 1 0 0 0
1 U
3835 0 0
2
45461.5 15
0
9 CA 7-Seg~
184 450 165 0 18 19
10 45 44 43 42 41 40 39 126 127
0 0 0 0 0 0 2 2 2
0
0 0 21104 0
7 AMBERCA
9 -41 58 -33
5 DISP3
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
3670 0 0
2
45461.5 16
0
6 74LS47
187 382 276 0 14 29
0 36 37 7 38 128 129 39 40 41
42 43 44 45 130
0
0 0 4848 0
6 74LS47
-21 -60 21 -52
2 U6
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
5616 0 0
2
45461.5 17
0
9 2-In AND~
219 823 314 0 3 22
0 55 54 4
0
0 0 624 180
6 74LS08
-21 -24 21 -16
3 U3B
-13 -25 8 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
9323 0 0
2
45461.5 18
0
6 74LS47
187 934 260 0 14 29
0 56 55 54 57 131 132 58 59 60
61 62 63 64 133
0
0 0 4848 0
6 74LS47
-21 -60 21 -52
2 U5
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
317 0 0
2
45461.5 19
0
9 CA 7-Seg~
184 1002 149 0 18 19
10 64 63 62 61 60 59 58 134 135
0 0 0 0 0 0 2 2 2
0
0 0 21104 0
7 AMBERCA
9 -41 58 -33
5 DISP2
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
3108 0 0
2
45461.5 20
0
7 74LS193
137 819 216 0 14 29
0 12 136 137 4 138 139 140 141 142
143 56 55 54 57
0
0 0 4848 0
7 74LS193
-24 -51 25 -43
2 U4
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
122 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 5 4 11 14 9 10 1 15 12
13 7 6 2 3 5 4 11 14 9
10 1 15 12 13 7 6 2 3 0
65 0 0 512 1 0 0 0
1 U
4299 0 0
2
45461.5 21
0
9 2-In AND~
219 1101 303 0 3 22
0 65 66 12
0
0 0 624 180
6 74LS08
-21 -24 21 -16
3 U3A
-13 -25 8 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
9672 0 0
2
45461.5 22
0
7 74LS193
137 1094 204 0 14 29
0 13 144 145 12 146 147 148 149 150
151 66 67 65 68
0
0 0 4848 0
7 74LS193
-24 -51 25 -43
2 U1
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
122 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 5 4 11 14 9 10 1 15 12
13 7 6 2 3 5 4 11 14 9
10 1 15 12 13 7 6 2 3 0
65 0 0 512 1 0 0 0
1 U
7876 0 0
2
45461.5 23
0
9 CA 7-Seg~
184 1277 137 0 18 19
10 75 74 73 72 71 70 69 152 153
0 0 0 0 0 0 2 2 2
0
0 0 21104 0
7 AMBERCA
9 -41 58 -33
5 DISP1
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
6369 0 0
2
45461.5 24
0
6 74LS47
187 1209 248 0 14 29
0 66 67 65 68 154 155 69 70 71
72 73 74 75 156
0
0 0 4848 0
6 74LS47
-21 -60 21 -52
2 U2
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
9172 0 0
2
45461.5 25
0
92
0 7 3 0 0 4096 0 0 1 36 0 3
1905 173
1905 163
1906 163
0 1 4 0 0 8320 0 0 14 65 0 8
777 313
699 313
699 191
584 191
584 142
496 142
496 193
510 193
0 1 5 0 0 4224 0 0 15 11 0 4
483 342
216 342
216 205
235 205
0 4 6 0 0 4224 0 0 15 7 0 4
474 425
221 425
221 232
235 232
0 1 7 0 0 4224 0 0 2 45 0 4
338 258
338 493
465 493
465 484
0 2 8 0 0 4224 0 0 2 55 0 4
620 237
620 493
483 493
483 484
1 3 6 0 0 0 0 3 2 0 0 2
474 405
474 439
2 3 9 0 0 8320 0 3 4 0 0 4
492 405
492 417
593 417
593 407
0 2 10 0 0 4224 0 0 4 56 0 2
584 247
584 362
0 1 11 0 0 4224 0 0 4 54 0 2
602 228
602 362
4 3 5 0 0 0 0 14 3 0 0 3
510 220
483 220
483 359
1 0 12 0 0 12416 0 21 0 0 79 6
787 189
768 189
768 334
1047 334
1047 303
1052 303
1 0 13 0 0 12416 0 23 0 0 15 6
1062 177
1040 177
1040 323
1385 323
1385 307
1390 307
0 1 14 0 0 12416 0 0 8 29 0 6
1665 299
1589 299
1589 353
1376 353
1376 185
1400 185
4 3 13 0 0 0 0 8 11 0 0 4
1400 212
1390 212
1390 310
1409 310
0 2 15 0 0 4224 0 0 11 20 0 3
1496 238
1496 301
1454 301
2 1 16 0 0 8320 0 10 11 0 0 4
1515 229
1503 229
1503 319
1454 319
1 11 17 0 0 4224 0 10 8 0 0 4
1515 220
1488 220
1488 221
1464 221
2 12 16 0 0 0 0 10 8 0 0 4
1515 229
1488 229
1488 230
1464 230
3 13 15 0 0 0 0 10 8 0 0 4
1515 238
1488 238
1488 239
1464 239
14 4 18 0 0 4224 0 8 10 0 0 4
1464 248
1507 248
1507 247
1515 247
7 7 19 0 0 4224 0 10 9 0 0 3
1585 220
1630 220
1630 181
8 6 20 0 0 8320 0 10 9 0 0 3
1585 229
1624 229
1624 181
9 5 21 0 0 8320 0 10 9 0 0 3
1585 238
1618 238
1618 181
10 4 22 0 0 8320 0 10 9 0 0 3
1585 247
1612 247
1612 181
11 3 23 0 0 8320 0 10 9 0 0 3
1585 256
1606 256
1606 181
12 2 24 0 0 8320 0 10 9 0 0 3
1585 265
1600 265
1600 181
1 13 25 0 0 4224 0 9 10 0 0 3
1594 181
1594 274
1585 274
4 3 14 0 0 0 0 6 7 0 0 4
1675 200
1665 200
1665 299
1687 299
0 1 26 0 0 4224 0 0 7 34 0 3
1776 226
1776 308
1732 308
0 2 27 0 0 4224 0 0 7 32 0 3
1782 208
1782 290
1732 290
1 11 27 0 0 0 0 5 6 0 0 4
1790 208
1763 208
1763 209
1739 209
2 12 28 0 0 4224 0 5 6 0 0 4
1790 217
1763 217
1763 218
1739 218
3 13 26 0 0 0 0 5 6 0 0 4
1790 226
1763 226
1763 227
1739 227
14 4 29 0 0 4224 0 6 5 0 0 4
1739 236
1782 236
1782 235
1790 235
7 0 3 0 0 4224 0 5 0 0 0 3
1860 208
1905 208
1905 169
8 6 30 0 0 8320 0 5 1 0 0 3
1860 217
1900 217
1900 163
9 5 31 0 0 8320 0 5 1 0 0 3
1860 226
1894 226
1894 163
10 4 32 0 0 8320 0 5 1 0 0 3
1860 235
1888 235
1888 163
11 3 33 0 0 8320 0 5 1 0 0 3
1860 244
1882 244
1882 163
12 2 34 0 0 8320 0 5 1 0 0 3
1860 253
1876 253
1876 163
1 13 35 0 0 4224 0 1 5 0 0 3
1870 163
1870 262
1860 262
1 11 36 0 0 4224 0 17 15 0 0 4
350 240
323 240
323 241
299 241
2 12 37 0 0 4224 0 17 15 0 0 4
350 249
323 249
323 250
299 250
3 13 7 0 0 0 0 17 15 0 0 4
350 258
323 258
323 259
299 259
14 4 38 0 0 4224 0 15 17 0 0 4
299 268
342 268
342 267
350 267
7 7 39 0 0 4224 0 17 16 0 0 3
420 240
465 240
465 201
8 6 40 0 0 8320 0 17 16 0 0 3
420 249
459 249
459 201
9 5 41 0 0 8320 0 17 16 0 0 3
420 258
453 258
453 201
10 4 42 0 0 8320 0 17 16 0 0 3
420 267
447 267
447 201
11 3 43 0 0 8320 0 17 16 0 0 3
420 276
441 276
441 201
12 2 44 0 0 8320 0 17 16 0 0 3
420 285
435 285
435 201
1 13 45 0 0 4224 0 16 17 0 0 3
429 201
429 294
420 294
1 11 11 0 0 0 0 12 14 0 0 4
625 228
598 228
598 229
574 229
2 12 8 0 0 0 0 12 14 0 0 4
625 237
598 237
598 238
574 238
3 13 10 0 0 0 0 12 14 0 0 4
625 246
598 246
598 247
574 247
14 4 46 0 0 4224 0 14 12 0 0 4
574 256
617 256
617 255
625 255
7 7 47 0 0 4224 0 12 13 0 0 3
695 228
740 228
740 189
8 6 48 0 0 8320 0 12 13 0 0 3
695 237
734 237
734 189
9 5 49 0 0 8320 0 12 13 0 0 3
695 246
728 246
728 189
10 4 50 0 0 8320 0 12 13 0 0 3
695 255
722 255
722 189
11 3 51 0 0 8320 0 12 13 0 0 3
695 264
716 264
716 189
12 2 52 0 0 8320 0 12 13 0 0 3
695 273
710 273
710 189
1 13 53 0 0 4224 0 13 12 0 0 3
704 189
704 282
695 282
4 3 4 0 0 0 0 21 18 0 0 4
787 216
777 216
777 314
796 314
0 2 54 0 0 4224 0 0 18 70 0 3
883 242
883 305
841 305
2 1 55 0 0 8320 0 19 18 0 0 4
902 233
890 233
890 323
841 323
1 11 56 0 0 4224 0 19 21 0 0 4
902 224
875 224
875 225
851 225
2 12 55 0 0 0 0 19 21 0 0 4
902 233
875 233
875 234
851 234
3 13 54 0 0 0 0 19 21 0 0 4
902 242
875 242
875 243
851 243
14 4 57 0 0 4224 0 21 19 0 0 4
851 252
894 252
894 251
902 251
7 7 58 0 0 4224 0 19 20 0 0 3
972 224
1017 224
1017 185
8 6 59 0 0 8320 0 19 20 0 0 3
972 233
1011 233
1011 185
9 5 60 0 0 8320 0 19 20 0 0 3
972 242
1005 242
1005 185
10 4 61 0 0 8320 0 19 20 0 0 3
972 251
999 251
999 185
11 3 62 0 0 8320 0 19 20 0 0 3
972 260
993 260
993 185
12 2 63 0 0 8320 0 19 20 0 0 3
972 269
987 269
987 185
1 13 64 0 0 4224 0 20 19 0 0 3
981 185
981 278
972 278
4 3 12 0 0 0 0 23 22 0 0 4
1062 204
1052 204
1052 303
1074 303
0 1 65 0 0 4224 0 0 22 84 0 3
1163 230
1163 312
1119 312
0 2 66 0 0 4224 0 0 22 82 0 3
1169 212
1169 294
1119 294
1 11 66 0 0 0 0 25 23 0 0 4
1177 212
1150 212
1150 213
1126 213
2 12 67 0 0 4224 0 25 23 0 0 4
1177 221
1150 221
1150 222
1126 222
3 13 65 0 0 0 0 25 23 0 0 4
1177 230
1150 230
1150 231
1126 231
14 4 68 0 0 4224 0 23 25 0 0 4
1126 240
1169 240
1169 239
1177 239
7 7 69 0 0 4224 0 25 24 0 0 3
1247 212
1292 212
1292 173
8 6 70 0 0 8320 0 25 24 0 0 3
1247 221
1286 221
1286 173
9 5 71 0 0 8320 0 25 24 0 0 3
1247 230
1280 230
1280 173
10 4 72 0 0 8320 0 25 24 0 0 3
1247 239
1274 239
1274 173
11 3 73 0 0 8320 0 25 24 0 0 3
1247 248
1268 248
1268 173
12 2 74 0 0 8320 0 25 24 0 0 3
1247 257
1262 257
1262 173
1 13 75 0 0 4224 0 24 25 0 0 3
1256 173
1256 266
1247 266
7
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 15
1199 50 1334 74
1206 55 1326 71
15 minutos(unidad)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 15
931 62 1066 86
938 67 1058 83
15 minutos(decena)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 13
647 66 766 90
654 71 758 87
13 horas(unidad)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 13
379 78 498 102
386 83 490 99
13 horas(decena)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 16
1546 17 1689 41
1553 22 1681 38
16 segundos(decena)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 16
1812 13 1955 37
1819 18 1947 34
16 segundos(unidad)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 18
996 3 1155 27
1003 8 1147 24
18 en cpu va la se�al
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
