CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 10 30 150 10
176 80 1438 831
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
43
13 Logic Switch~
5 64 179 0 10 11
0 7 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V8
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
5.90124e-315 0
0
13 Logic Switch~
5 64 137 0 1 11
0 8
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V7
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
391 0 0
2
5.90124e-315 5.26354e-315
0
13 Logic Switch~
5 63 94 0 1 11
0 9
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V6
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3124 0 0
2
5.90124e-315 5.30499e-315
0
13 Logic Switch~
5 65 49 0 1 11
0 10
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3421 0 0
2
5.90124e-315 5.32571e-315
0
13 Logic Switch~
5 88 234 0 10 11
0 3 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
8157 0 0
2
5.90124e-315 5.34643e-315
0
13 Logic Switch~
5 88 443 0 1 11
0 6
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5572 0 0
2
5.90124e-315 5.3568e-315
0
13 Logic Switch~
5 92 362 0 1 11
0 5
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8901 0 0
2
5.90124e-315 5.36716e-315
0
13 Logic Switch~
5 94 294 0 10 11
0 4 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
7361 0 0
2
5.90124e-315 5.37752e-315
0
7 Ground~
168 129 741 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4747 0 0
2
45434.5 0
0
9 CA 7-Seg~
184 387 651 0 18 19
10 17 16 15 14 13 12 11 40 41
0 0 0 0 2 2 0 2 2
0
0 0 21088 0
5 REDCA
16 -41 51 -33
5 DISP2
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
972 0 0
2
45434.5 1
0
9 CA 7-Seg~
184 384 510 0 18 19
10 24 23 22 21 20 19 18 42 43
0 0 0 0 0 0 0 2 2
0
0 0 21088 0
5 REDCA
16 -41 51 -33
5 DISP1
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
3472 0 0
2
45434.5 2
0
6 74LS47
187 214 676 0 14 29
0 6 5 4 3 44 2 11 12 13
14 15 16 17 25
0
0 0 4848 0
6 74LS47
-21 -60 21 -52
2 U6
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
9998 0 0
2
5.90124e-315 5.38788e-315
0
6 74LS47
187 209 527 0 14 29
0 7 8 9 10 45 25 18 19 20
21 22 23 24 46
0
0 0 4848 0
6 74LS47
-21 -60 21 -52
2 U5
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
3536 0 0
2
5.90124e-315 5.39306e-315
0
14 Logic Display~
6 694 53 0 1 2
10 26
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L16
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4597 0 0
2
45434.5 3
0
14 Logic Display~
6 691 108 0 1 2
10 27
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L15
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3835 0 0
2
45434.5 4
0
14 Logic Display~
6 690 160 0 1 2
10 28
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L14
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3670 0 0
2
45434.5 5
0
9 2-In XOR~
219 530 63 0 3 22
0 30 27 26
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U4C
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 5 0
1 U
5616 0 0
2
45434.5 6
0
9 2-In XOR~
219 528 130 0 3 22
0 31 28 27
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U4B
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 5 0
1 U
9323 0 0
2
45434.5 7
0
9 2-In XOR~
219 528 186 0 3 22
0 32 29 28
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U4A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 5 0
1 U
317 0 0
2
45434.5 8
0
14 Logic Display~
6 705 218 0 1 2
10 29
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L13
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3108 0 0
2
45434.5 9
0
9 2-In XOR~
219 526 256 0 3 22
0 33 34 29
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U3D
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 4 0
1 U
4299 0 0
2
45434.5 10
0
9 2-In XOR~
219 522 323 0 3 22
0 35 36 34
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U3C
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 4 0
1 U
9672 0 0
2
45434.5 11
0
14 Logic Display~
6 699 272 0 1 2
10 34
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L12
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7876 0 0
2
45434.5 12
0
9 2-In XOR~
219 520 374 0 3 22
0 37 38 36
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U3B
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 4 0
1 U
6369 0 0
2
45434.5 13
0
14 Logic Display~
6 701 310 0 1 2
10 36
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L11
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9172 0 0
2
45434.5 14
0
14 Logic Display~
6 702 360 0 1 2
10 38
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L10
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7100 0 0
2
45434.5 15
0
9 2-In XOR~
219 521 418 0 3 22
0 39 6 38
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U3A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
3820 0 0
2
45434.5 16
0
14 Logic Display~
6 643 421 0 1 2
10 6
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L9
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7678 0 0
2
45434.5 17
0
14 Logic Display~
6 450 240 0 1 2
10 35
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
961 0 0
2
5.90124e-315 5.39824e-315
0
9 2-In XOR~
219 317 283 0 3 22
0 3 4 35
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U1D
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 3 0
1 U
3178 0 0
2
5.90124e-315 5.40342e-315
0
14 Logic Display~
6 448 413 0 1 2
10 6
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L8
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3409 0 0
2
5.90124e-315 5.4086e-315
0
14 Logic Display~
6 450 355 0 1 2
10 39
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L7
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3951 0 0
2
5.90124e-315 5.41378e-315
0
9 2-In XOR~
219 277 391 0 3 22
0 5 6 39
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U1C
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 3 0
1 U
8885 0 0
2
5.90124e-315 5.41896e-315
0
14 Logic Display~
6 449 305 0 1 2
10 37
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3780 0 0
2
5.90124e-315 5.42414e-315
0
9 2-In XOR~
219 279 334 0 3 22
0 4 5 37
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U1B
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
9265 0 0
2
5.90124e-315 5.42933e-315
0
14 Logic Display~
6 449 194 0 1 2
10 33
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9442 0 0
2
5.90124e-315 5.43192e-315
0
9 2-In XOR~
219 275 220 0 3 22
0 7 3 33
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U2D
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 2 0
1 U
9424 0 0
2
5.90124e-315 5.43451e-315
0
9 2-In XOR~
219 276 169 0 3 22
0 8 7 32
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U2C
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 2 0
1 U
9968 0 0
2
5.90124e-315 5.4371e-315
0
14 Logic Display~
6 449 145 0 1 2
10 32
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9281 0 0
2
5.90124e-315 5.43969e-315
0
14 Logic Display~
6 447 99 0 1 2
10 31
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8464 0 0
2
5.90124e-315 5.44228e-315
0
9 2-In XOR~
219 277 120 0 3 22
0 9 8 31
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U2B
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
7168 0 0
2
5.90124e-315 5.44487e-315
0
14 Logic Display~
6 447 47 0 1 2
10 30
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3171 0 0
2
5.90124e-315 5.44746e-315
0
9 2-In XOR~
219 272 70 0 3 22
0 10 9 30
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U2A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
4139 0 0
2
5.90124e-315 5.45005e-315
0
69
6 1 2 0 0 4224 0 12 9 0 0 3
182 721
129 721
129 735
0 4 3 0 0 4224 0 0 12 59 0 3
114 234
114 667
182 667
0 3 4 0 0 4224 0 0 12 56 0 3
126 294
126 658
182 658
0 2 5 0 0 8320 0 0 12 54 0 4
113 361
152 361
152 649
182 649
0 1 6 0 0 4224 0 0 12 51 0 3
147 443
147 640
182 640
0 1 7 0 0 4224 0 0 13 62 0 5
177 169
177 472
164 472
164 491
177 491
0 2 8 0 0 4224 0 0 13 65 0 3
155 133
155 500
177 500
0 3 9 0 0 4224 0 0 13 68 0 3
137 89
137 509
177 509
0 4 10 0 0 4224 0 0 13 69 0 3
169 53
169 518
177 518
7 7 11 0 0 8320 0 12 10 0 0 5
252 640
331 640
331 723
402 723
402 687
8 6 12 0 0 4224 0 12 10 0 0 5
252 649
336 649
336 718
396 718
396 687
9 5 13 0 0 4224 0 12 10 0 0 5
252 658
341 658
341 713
390 713
390 687
10 4 14 0 0 4224 0 12 10 0 0 5
252 667
346 667
346 708
384 708
384 687
11 3 15 0 0 4224 0 12 10 0 0 5
252 676
351 676
351 703
378 703
378 687
12 2 16 0 0 4224 0 12 10 0 0 5
252 685
356 685
356 698
372 698
372 687
13 1 17 0 0 4224 0 12 10 0 0 3
252 694
366 694
366 687
7 7 18 0 0 8320 0 13 11 0 0 5
247 491
324 491
324 584
399 584
399 546
8 6 19 0 0 4224 0 13 11 0 0 5
247 500
329 500
329 579
393 579
393 546
9 5 20 0 0 4224 0 13 11 0 0 5
247 509
334 509
334 574
387 574
387 546
10 4 21 0 0 4224 0 13 11 0 0 5
247 518
339 518
339 569
381 569
381 546
11 3 22 0 0 4224 0 13 11 0 0 5
247 527
344 527
344 564
375 564
375 546
12 2 23 0 0 4224 0 13 11 0 0 5
247 536
349 536
349 559
369 559
369 546
13 1 24 0 0 4224 0 13 11 0 0 5
247 545
354 545
354 554
363 554
363 546
6 14 25 0 0 8320 0 13 12 0 0 6
177 572
173 572
173 736
260 736
260 721
246 721
3 1 26 0 0 8320 0 17 14 0 0 4
563 63
563 69
694 69
694 71
0 2 27 0 0 8320 0 0 17 27 0 5
600 130
600 83
506 83
506 72
514 72
3 1 27 0 0 0 0 18 15 0 0 5
561 130
652 130
652 108
691 108
691 126
0 2 28 0 0 8192 0 0 18 29 0 5
588 186
588 150
504 150
504 139
512 139
3 1 28 0 0 4224 0 19 16 0 0 5
561 186
650 186
650 184
690 184
690 178
0 2 29 0 0 8192 0 0 19 34 0 5
586 256
586 206
504 206
504 195
512 195
1 1 30 0 0 4096 0 17 42 0 0 5
514 54
459 54
459 73
447 73
447 65
1 1 31 0 0 8192 0 40 18 0 0 3
447 117
447 121
512 121
1 1 32 0 0 8192 0 39 19 0 0 3
449 163
449 177
512 177
3 1 29 0 0 4224 0 21 20 0 0 6
559 256
649 256
649 235
667 235
667 236
705 236
1 1 33 0 0 8192 0 36 21 0 0 5
449 212
449 225
502 225
502 247
510 247
0 2 34 0 0 4224 0 0 21 37 0 4
609 276
497 276
497 265
510 265
3 1 34 0 0 0 0 22 23 0 0 6
555 323
609 323
609 253
622 253
622 290
699 290
0 1 35 0 0 4096 0 0 22 48 0 4
450 268
500 268
500 314
506 314
2 0 36 0 0 12416 0 22 0 0 40 5
506 332
504 332
504 323
591 323
591 298
3 1 36 0 0 0 0 24 25 0 0 8
553 374
591 374
591 298
604 298
604 310
651 310
651 328
701 328
0 1 37 0 0 8192 0 0 24 53 0 5
448 334
448 327
494 327
494 365
504 365
0 2 38 0 0 8192 0 0 24 43 0 4
572 374
572 316
504 316
504 383
1 3 38 0 0 8320 0 26 27 0 0 5
702 378
702 374
572 374
572 418
554 418
2 0 6 0 0 0 0 27 0 0 46 3
505 427
493 427
493 440
1 0 39 0 0 4096 0 27 0 0 50 4
505 409
462 409
462 376
450 376
1 1 6 0 0 0 0 31 28 0 0 4
448 431
448 440
643 440
643 439
0 1 9 0 0 0 0 0 3 68 0 3
105 89
105 94
75 94
3 1 35 0 0 4224 0 30 29 0 0 3
350 283
450 283
450 258
0 1 6 0 0 0 0 0 31 51 0 3
253 434
448 434
448 431
3 1 39 0 0 4224 0 33 32 0 0 3
310 391
450 391
450 373
1 2 6 0 0 0 0 6 33 0 0 4
100 443
253 443
253 400
261 400
0 1 5 0 0 0 0 0 33 54 0 3
210 343
210 382
261 382
3 1 37 0 0 4224 0 35 34 0 0 3
312 334
449 334
449 323
2 1 5 0 0 0 0 35 7 0 0 4
263 343
113 343
113 362
104 362
0 1 4 0 0 0 0 0 35 56 0 3
232 294
232 325
263 325
1 2 4 0 0 0 0 8 30 0 0 4
106 294
262 294
262 292
301 292
0 1 3 0 0 0 0 0 30 59 0 5
237 231
237 276
262 276
262 274
301 274
3 1 33 0 0 4224 0 37 36 0 0 3
308 220
449 220
449 212
1 2 3 0 0 0 0 5 37 0 0 6
100 234
115 234
115 231
251 231
251 229
259 229
0 1 7 0 0 0 0 0 37 62 0 3
186 169
186 211
259 211
3 1 32 0 0 4224 0 38 39 0 0 3
309 169
449 169
449 163
1 2 7 0 0 0 0 1 38 0 0 6
76 179
107 179
107 169
252 169
252 178
260 178
0 1 8 0 0 0 0 0 38 65 0 3
229 133
229 160
260 160
3 1 31 0 0 4224 0 41 40 0 0 3
310 120
447 120
447 117
1 2 8 0 0 0 0 2 41 0 0 6
76 137
106 137
106 133
253 133
253 129
261 129
0 1 9 0 0 0 0 0 41 68 0 3
193 89
193 111
261 111
3 1 30 0 0 4224 0 43 42 0 0 3
305 70
447 70
447 65
0 2 9 0 0 0 0 0 43 0 0 4
101 89
202 89
202 79
256 79
1 1 10 0 0 0 0 4 43 0 0 6
77 49
95 49
95 53
202 53
202 61
256 61
12
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 12
571 -4 688 20
581 4 677 20
12 gray-binario
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
26 38 55 62
36 46 44 62
1 A
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
26 75 55 99
36 83 44 99
1 B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
27 119 56 143
37 127 45 143
1 C
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
27 155 56 179
37 163 45 179
1 D
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
30 217 59 241
40 225 48 241
1 E
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
35 279 64 303
45 287 53 303
1 F
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
39 341 68 365
49 349 57 365
1 G
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
31 426 60 450
41 434 49 450
1 H
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 12
202 -3 319 21
212 5 308 21
12 binario-gray
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 22
116 774 307 798
123 779 299 795
22 BCD a display de 7 seg
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 14
145 796 272 820
152 802 264 818
14 decodificacion
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
