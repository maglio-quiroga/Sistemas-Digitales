CircuitMaker Text
5.6
Probes: 1
c4[p]
Transient Analysis
0 989 286 65280
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 90 30 110 10
176 80 1534 795
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
176 80 1534 437
9961490 0
0
6 Title:
5 Name:
0
0
0
22
10 555 Timer~
219 936 233 0 8 17
0 2 5 4 3 6 7 7 3
0
0 0 4944 0
3 555
-11 -36 10 -28
2 U2
-7 -46 7 -38
0
0
29 %D %1 %2 %3 %4 %5 %6 %7 %8 %S
0
0
4 DIP8
17

0 1 2 3 4 5 6 7 8 1
2 3 4 5 6 7 8 0
88 0 0 0 1 0 0 0
1 U
3284 0 0
2
45450.7 10
0
2 +V
167 1013 112 0 1 3
0 3
0
0 0 54256 0
2 5V
-8 -21 6 -13
2 V4
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
659 0 0
2
45450.7 9
0
10 Capacitor~
219 985 285 0 2 5
0 2 7
0
0 0 848 90
3 9uF
12 -1 33 7
2 C4
13 -8 27 0
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
3800 0 0
2
45450.7 8
0
7 Ground~
168 985 325 0 1 3
0 2
0
0 0 53360 0
0
5 GND10
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6792 0 0
2
45450.7 7
0
7 Ground~
168 1047 327 0 1 3
0 2
0
0 0 53360 0
0
4 GND9
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3701 0 0
2
45450.7 6
0
10 Capacitor~
219 1047 287 0 2 5
0 2 6
0
0 0 848 90
6 0.01uF
1 0 43 8
2 C3
15 -10 29 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
6316 0 0
2
45450.7 5
0
7 Ground~
168 787 195 0 1 3
0 2
0
0 0 53360 270
0
4 GND8
-14 -28 14 -20
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8734 0 0
2
45450.7 4
0
11 Signal Gen~
195 690 303 0 64 64
0 5 2 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1092616192 0 1084227584
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 266
20
1 10 0 5 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
5 -5/5V
-18 -30 17 -22
2 V2
-7 -40 7 -32
0
0
36 %D %1 %2 DC 0 SIN(0 5 10 0 0) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 0 0 0 0
1 V
7988 0 0
2
45450.7 3
0
7 Ground~
168 740 354 0 1 3
0 2
0
0 0 53360 0
0
4 GND7
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
3217 0 0
2
45450.7 2
0
4 LED~
171 747 216 0 2 2
10 4 2
0
0 0 880 180
4 LED1
16 0 44 8
2 D2
23 -10 37 -2
0
0
11 %D %1 %2 %M
0
0
0
5

0 1 2 1 2 0
68 0 0 0 0 0 0 0
1 D
3965 0 0
2
45450.7 1
0
4 LED~
171 282 245 0 2 2
10 9 2
0
0 0 880 180
4 LED1
16 0 44 8
2 D1
23 -10 37 -2
0
0
11 %D %1 %2 %M
0
0
0
5

0 1 2 1 2 0
68 0 0 0 0 0 0 0
1 D
8239 0 0
2
45450.7 0
0
7 Ground~
168 275 383 0 1 3
0 2
0
0 0 53360 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
828 0 0
2
45450.7 0
0
11 Signal Gen~
195 225 332 0 19 64
0 10 2 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1092616192 0 1084227584
20
1 10 0 5 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
5 -5/5V
-18 -30 17 -22
2 V3
-7 -40 7 -32
0
0
36 %D %1 %2 DC 0 SIN(0 5 10 0 0) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 0 0 0 0
1 V
6187 0 0
2
45450.7 0
0
7 Ground~
168 322 224 0 1 3
0 2
0
0 0 53360 270
0
4 GND3
-14 -28 14 -20
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7107 0 0
2
5.90126e-315 0
0
10 Capacitor~
219 582 316 0 2 5
0 2 11
0
0 0 848 90
6 0.01uF
1 0 43 8
2 C2
15 -10 29 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
6433 0 0
2
5.90126e-315 5.26354e-315
0
7 Ground~
168 582 356 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8559 0 0
2
5.90126e-315 0
0
7 Ground~
168 520 354 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3674 0 0
2
5.90126e-315 0
0
10 Capacitor~
219 520 314 0 2 5
0 2 12
0
0 0 848 90
5 4.5uF
5 -1 40 7
2 C1
13 -8 27 0
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
5697 0 0
2
5.90126e-315 0
0
2 +V
167 548 141 0 1 3
0 8
0
0 0 54256 0
2 5V
-8 -21 6 -13
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3805 0 0
2
5.90126e-315 0
0
10 555 Timer~
219 471 262 0 8 17
0 2 10 9 8 11 12 12 8
0
0 0 4944 0
3 555
-11 -36 10 -28
2 U1
-7 -46 7 -38
0
0
29 %D %1 %2 %3 %4 %5 %6 %7 %8 %S
0
0
4 DIP8
17

0 1 2 3 4 5 6 7 8 1
2 3 4 5 6 7 8 0
88 0 0 0 1 0 0 0
1 U
5219 0 0
2
5.90126e-315 0
0
9 Resistor~
219 985 182 0 4 5
0 7 3 0 1
0
0 0 880 90
2 2k
9 -1 23 7
2 R2
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3795 0 0
2
45450.7 11
0
9 Resistor~
219 520 211 0 4 5
0 12 8 0 1
0
0 0 880 90
2 1k
9 -1 23 7
2 R1
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3637 0 0
2
5.90126e-315 0
0
28
2 0 2 0 0 8192 0 10 0 0 7 4
749 206
749 167
843 167
843 196
2 0 2 0 0 8320 0 11 0 0 20 4
284 235
284 170
379 170
379 225
4 0 3 0 0 8208 0 1 0 0 13 4
904 251
887 251
887 151
985 151
3 1 4 0 0 4240 0 1 10 0 0 3
904 242
749 242
749 226
1 2 2 0 0 16 0 9 8 0 0 3
740 348
740 308
721 308
2 1 5 0 0 12432 0 1 8 0 0 4
904 233
820 233
820 298
721 298
1 1 2 0 0 144 0 1 7 0 0 4
904 224
855 224
855 196
794 196
5 2 6 0 0 4240 0 1 6 0 0 3
968 251
1047 251
1047 278
1 1 2 0 0 16 0 6 5 0 0 2
1047 296
1047 321
1 1 2 0 0 16 0 3 4 0 0 2
985 294
985 319
6 0 7 0 0 4112 0 1 0 0 12 2
968 242
985 242
0 2 7 0 0 4240 0 0 3 14 0 2
985 233
985 276
2 0 3 0 0 16 0 21 0 0 15 3
985 164
985 151
1013 151
7 1 7 0 0 16 0 1 21 0 0 3
968 233
985 233
985 200
8 1 3 0 0 8336 0 1 2 0 0 3
968 224
1013 224
1013 121
4 0 8 0 0 8192 0 20 0 0 26 4
439 280
422 280
422 180
520 180
3 1 9 0 0 4224 0 20 11 0 0 3
439 271
284 271
284 255
1 2 2 0 0 0 0 12 13 0 0 3
275 377
275 337
256 337
2 1 10 0 0 12416 0 20 13 0 0 4
439 262
355 262
355 327
256 327
1 1 2 0 0 128 0 20 14 0 0 4
439 253
390 253
390 225
329 225
5 2 11 0 0 4224 0 20 15 0 0 3
503 280
582 280
582 307
1 1 2 0 0 0 0 15 16 0 0 2
582 325
582 350
1 1 2 0 0 0 0 18 17 0 0 2
520 323
520 348
6 0 12 0 0 4096 0 20 0 0 25 2
503 271
520 271
0 2 12 0 0 4224 0 0 18 27 0 2
520 262
520 305
2 0 8 0 0 0 0 22 0 0 28 3
520 193
520 180
548 180
7 1 12 0 0 0 0 20 22 0 0 3
503 262
520 262
520 229
8 1 8 0 0 8320 0 20 19 0 0 3
503 253
548 253
548 150
1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 22
104 74 299 96
113 81 289 97
22 Temps 555 monoestables
0
2065 0 1
0
0
2 V1
1 0 -1
0
0 0 0
3 0 1 4
0 0.5 0.002 0.002
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
14112 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
